module i2c_write_tb();

    reg         rst_n       ;
    reg         clk         ;
    reg         pre_ready   ;
    reg [7:0]   pre_data    ;
    reg [6:0]   i2c_slave_addr;
    wire        i2c_busy    ;
    wire        











endmodule

